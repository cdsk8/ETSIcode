��  CCircuit��  CSerializeHack           ��  CPart              ���  CEarth�� 	 CTerminal  p@�A                �NJ)f?    �4�L        ��      �
�  4 HI I                �NJ)f�    , :4 R        ��      �� 	 CResistor��  CValue  (    1800         �@      �?   
�  $9                �4r�+Jb�  
�  �        -`��0@�4r�+Jb?    $        ��      ��  0^Pl    6800        ��@      �?   
�  Lpaq                ���f�>�  
�   p5q        �bg�k	@���f�>?    4lLt        ��      ��  �^ l    1800         �@      �?   
�  �pq        �bg�k	@���f�>�  
�  �p�q        -`��0@���f�>?    �l�t        ��      ��   ^ l    8200        �@      �?   
�  p1q        -`��0@?Cp��U�  
�  � pq             .@?Cp��U?    lt        ��      ��  Pp    5600        �@      �?   
�  l�        -`��0@��Y$gKV�  
�  @U       �$��#G'@��Y$gKV?    Tl    "    ��      ��        270        �p@      �?   
�  1       �$��#G'@��Y$gKV�  
�  �        N��@(@��Y$gKV?        &    ��      ��  � �     2200        0�@      �?   
�  � �        N��@(@��Y$gKV�  
�  � �              .@��Y$gKV?    � �     *    ��      ��  CBattery�  T /| =    15V         .@      �? V 
�  t H� I             .@�NJ)f�  
�  H H] I      	         �NJ)f?    \ <t T    /    ��                    ���  CWire  pqA       2�  p@qq       2�  �@�q       2�  ��A       2�  �@�A      2�  ��A       2�  �@�q       2�  p!q      2�  `pqq      2�  8q      2�  �p�q      2�  ��      2�  ��      2�  0p�q      2�  0A      2�  � �       2�  � p� q      2�  � H� q       2�  � �       2�  � � I                     �                             4    0   <  >    ;  :    :  =    @  C  " " ? # A # & & A ' B ' * * B + E + / / D 0  0 <  3 ; 6 = > 7 9 5 ? 7 8 @    4  3 5  6  " 8  9 & # * ' D  F C F + E /             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 