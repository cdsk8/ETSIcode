----------------------------------------------------------------------------------------------------------
--                              CIRCUITO ANTIRREBOTES POR RETARDO                              
----------------------------------------------------------------------------------------------------------
-- ESTE CIRCUITO ELIMINA LOS REBOTES MEDIANTE LA GENERACI�N DE RETARDOS.
-- PRODUCE UN �NICO FLANCO DE SUBIDA CADA VEZ QUE SE PRESIONA EL "PULSADOR". 
-- MODO DE CONEXI�N:
--   CLK_50MHZ: AL GENERADOR DE RELOJ DE 50 MHZ DE LA TARJETA (C9).
--   E: A UNO DE LOS PULSADORES SIGUIENTES DE LA TARJETA:
--       BTN CENTER (K17).
--       BTN NORTH (V4).
--       BTN EAST (H13).
--       BTN SOUTH (K17).
--       BTN WEST (D18).
--   S: A LAS ENTRADAS DEL CIRCUITO QUE NECESITEN UNA SE�AL SIN REBOTES.

-- EN EL FICHERO DE RESTRICCIONES ".UCF" SE DEBEN A�ADIR LAS SENTENCIAS SIGUIENTES:
-- NET "CLK_50MHZ" LOC = C9;
-- NET "PULSADOR" LOC = "REFERENCIA DEL PULSADOR" | PULLDOWN;
-- NET "PULSADOR" CLOCK_DEDICATED_ROUTE = FALSE;

-- PARA SIMULAR EL SISTEMA DONDE SE INSERTE ESTE CIRCUITO, ASIGNAR AL PAR�METRO
-- "SIMULAR" DE GENERIC EL VALOR '1' ANTES DE SINTETIZAR.
-- PARA IMPLEMENTAR EN LA FPGA EL SISTEMA DONDE SE INSERTE ESTE CIRCUITO, ASIGNAR
-- AL PAR�METRO "SIMULAR" DE GENERIC EL VALOR '0' ANTES DE SINTETIZAR.
----------------------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ANTIRREBOTES IS
	GENERIC (SIMULAR: STD_LOGIC := '1');	--Cambiame cuando vallas a compilar
	PORT (CLK_50MHZ, E: IN STD_LOGIC; S: OUT STD_LOGIC);
END ANTIRREBOTES;

ARCHITECTURE A_ANTIRREBOTES OF ANTIRREBOTES IS

SIGNAL HC_1, HC_2, FC_1, FC_2: STD_LOGIC := '0';
SIGNAL CONTADOR_1, CONTADOR_2: STD_LOGIC_VECTOR (20 DOWNTO 0) := (OTHERS => '0');

BEGIN

WITH SIMULAR SELECT S <= E WHEN '1', HC_1 WHEN OTHERS;

PROCESS (FC_2, E)
BEGIN
	IF FC_2 = '1' THEN HC_1 <= '0';
	ELSIF E'EVENT AND E = '1' THEN HC_1 <= '1';
	END IF;
END PROCESS;

PROCESS (HC_1, CLK_50MHZ)
BEGIN
	IF HC_1 = '0' THEN CONTADOR_1 <= (OTHERS => '0');
	ELSIF FC_1 = '0' AND CLK_50MHZ'EVENT AND CLK_50MHZ = '1'
			THEN CONTADOR_1 <= CONTADOR_1 + 1;
	END IF;
END PROCESS;

FC_1 <= CONTADOR_1(20);	

PROCESS (FC_1, E)
BEGIN
	IF FC_1 = '0' THEN HC_2 <= '0';
	ELSIF E'EVENT AND E = '0' THEN HC_2 <= '1';
	END IF;
END PROCESS;
	
PROCESS (FC_1, CLK_50MHZ)
BEGIN
	IF FC_1 = '0' THEN CONTADOR_2 <= (OTHERS => '0');
	ELSIF HC_2 = '1' AND CLK_50MHZ'EVENT AND CLK_50MHZ = '1'
			THEN CONTADOR_2 <= CONTADOR_2 + 1;
	END IF;
END PROCESS;

FC_2 <= CONTADOR_2(20);
	
END A_ANTIRREBOTES;
