��  CCircuit��  CSerializeHack           ��  CPart    0   0     ��� 	 CResistor��  CValue  �n�|    680        @�@      �?   �� 	 CTerminal  ����        !�|��@�E(Bq?  �  ����     	       LI*>�E(Bq�    �|��        ��      �
�  �Y�g    100           Y@      �?   �  �@�U      
 	 �J�Y�J
@�E(Bq?  �  �l��      	 !�|��@�E(Bq�    �T�l         ��      �
�  �.�<    1k        @�@      �?k  �  �@�A     
   �J�Y�J
@�E(Bq�  �  �@�A        ��4   @�E(Bq?    �<�D        ��      ��  CBattery
�  kY�g    7.5V(          @      �? V �  �@�U       	 ��4   @�E(Bq�  �  �l��     	      LI*>�E(Bq?    �T�l         ��      �
�  � Yg    15V(          .@      �? V �  @U       	       .@�E(B��  �  l�                �E(B�?    T$l         ��      �
�  (.H<    1k        @�@      �?k  �  D@YA        e%+Y�J@�E(B��  �  @-A             .@�E(B�?    ,<DD    "    ��      �
�  3YSg    100           Y@      �?   �  X@YU       	 e%+Y�J@�E(B�?  �  XlY�      	 �u�{��@�E(B��    TT\l     &    ��      �
�  (nH|    680        @�@      �?   �  D�Y�        �u�{��@�E(B�?  �  �-�                 �E(B��    ,|D�    *    ��      �
�  � f� t    680        @�@      �?   �  � x� y       ��Ngm��~����i��  �  x x� y        �tQ�ԯ�?~����i�?    � t� |    .    ��      �
�  � Q� _    100           Y@      �?   �  � 8� M       	 j �f�~����i��  �  � d� y      	 ��Ngm��~����i�?    � L� d     2    ��      �
�  � &� 4    1k        @�@      �?k  �  � 8� 9       j �f�}����i�?  �  x 8� 9       I�K�"�(�}����i��    � 4� <    6    ��      ��  CVPulse�� 
 CSineValue  3 Qk _    1Hz8          �?      �? Hz       .@      �?                      �  x 8y M       	 I�K�"�(�����i�?  �  x dy y      	 �tQ�ԯ�?~����i��    l L� d     <    ��            0   0     �    0   0     �    0   0         0   0                              #    + " " & #  # & " & ' ' * * * ' +  + . . 3 / = / 2 6 2 3 3 . 6 6 2 7 < 7 < 7 < = = /           �5s�        @     +        @            4@    "V  (      �P                
         .@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 